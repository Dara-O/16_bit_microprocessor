`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/12/2021 08:39:56 PM
// Design Name: 
// Module Name: FSMStateDataPackage
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package FSMStateData; 
    
    typedef enum logic [3:0] {S0, S1, S2, S3, S4, S5, 
                              S6, S7, S8, S9, S10, S11} state_t;
                          
endpackage
